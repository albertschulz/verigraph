module parent();
    a i_a();
endmodule