module a();
endmodule;

module b();
endmodule;

module parent();

    a i_a();
    b i_a();

endmodule