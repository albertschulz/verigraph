package pkg;
endpackage

module parent();
    import pkg::*;
endmodule