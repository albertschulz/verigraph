interface intf;
endinterface

module a();
    intf i_intf();
endmodule